package mem_model_pkg;

    import uvm_pkg::*;
  
    `include "uvm_macros.svh"
    `include "mem_model.sv"
  
  endpackage