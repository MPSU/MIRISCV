`include "miriscv_riscv_instr_base_test.sv"
`include "miriscv_asm_program_gen.sv"
