//////////////////////////////////////
// Miriscv core environment package //
//////////////////////////////////////

package miriscv_test_pkg;

  import uvm_pkg::*;
  import miriscv_env_pkg::*;
  import miriscv_mem_intf_agent_pkg::*;
  import riscv_signature_pkg::*;

  `include "miriscv_report_server.sv"
  `include "miriscv_vseq.sv"
  `include "miriscv_base_test.sv"
  `include "miriscv_self_check_test_lib.sv"

endpackage