//////////////////////////////////////
// Miriscv core environment package //
//////////////////////////////////////

package miriscv_env_pkg;

  import uvm_pkg::*;
  import miriscv_mem_intf_agent_pkg::*;

  `include "miriscv_vseqr.sv"
  `include "miriscv_env.sv"

endpackage
