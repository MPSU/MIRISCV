/***********************************************************************************
 * Copyright (C) 2023 National Research University of Electronic Technology (MIET),
 * Institute of Microdevices and Control Systems.
 * See LICENSE file for licensing details.
 *
 * This file is a part of miriscv core.
 *
 ***********************************************************************************/

package  miriscv_cu_pkg;

  parameter NO_BYPASS = 2'd0;
  parameter BYPASS_E  = 2'd1;
  parameter BYPASS_M  = 2'd2;

endpackage :  miriscv_cu_pkg
